module andgate (a, b, y);
    input  a , b;
    output y;
    y = a & b;  
endmodule